`timescale 1ns / 1ps

module elem_eng(
	// TODO
);
	// TODO
endmodule
