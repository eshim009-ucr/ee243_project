`timescale 1ns / 1ps

module conv_eng(
	// TODO
);
	// TODO
endmodule
