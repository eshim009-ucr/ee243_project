`timescale 1ns / 1ps

module dpu(
	// TODO
);
	// TODO
endmodule
