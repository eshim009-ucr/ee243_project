`timescale 1ns / 1ps

module dwcv_eng(
	// TODO
);
	// TODO
endmodule
