`timescale 1ns / 1ps

module pool_eng(
	// TODO
);
	// TODO
endmodule
